reg q;
always @*
  q = sel ? a : b;
